module instr(addr, com);
    input [31:0] addr;
    output wire [31:0] com;
    reg [31:0] instr[31:0]; 
    initial begin
        instr[0] = 32'b100011_00000_00000_0000_0000_0000_0000;  // $0 = $0
        instr[1] = 32'b100011_00000_00001_0000_0000_0000_0001;  // $1 = $0 
        instr[2] = 32'b001000_00000_00000_0000_0000_0000_0001;  // $0 = $0 + 1;
        instr[3] = 32'b001000_00001_00001_0000_0000_0000_0011;  // $1 = $1 + 3
        instr[4] = 32'b001000_00000_00000_0000_0000_0000_0001;  // $0 = $0 + 1
        instr[5] = 32'b000000_00000_00001_00000_xxxxx_101010;   // $0 = ($0 == $1)
        instr[6] = 32'b000100_00000_00000_0000_0000_0000_0001;  // $0 == 0 
        instr[7] = 32'b001000_00001_00001_0000_0000_0000_1010;  // $1 = $1 + 5
        instr[8] = 32'b001000_00000_00000_0000_0000_0000_1010;  // $0 = $0 + 5
        instr[9] = 32'b101011_00011_00000_0000_0000_0000_0000;
    end
    assign com = instr[addr];
    
endmodule
